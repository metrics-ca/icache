`include "uvm_macros.svh"

package tb_icache_pkg;
import uvm_pkg::*;

`include "ic_xact.svh"

endpackage

