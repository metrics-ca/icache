`include "uvm_macros.svh"

package tb_dram_ctrl_pkg;
import uvm_pkg::*;

`include "dram_ctrl_xact.svh"
`include "dram_ctrl_monitor.svh"

endpackage